module display(clk,rst,innum,SEG0,SEG1);

input clk;
input rst;
input [5:0] innum;

output [6:0] SEG0;
output [6:0] SEG1;

reg [6:0] SEG0;
reg [6:0] SEG1;


endmodule